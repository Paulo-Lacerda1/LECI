library IEEE;
use IEEE.STD_LOGIC_1164.all;


entity name1 is
	
	port (wren, clk : in  std_logic;
		  dataIn    : in  std_logic_vector(7 downto 0);
		  dataOut   :   out std_logic_vector(7 downto 0));
	
end name1;

architecture Behavioral of name1 is
begin

	process(clk)
	
	begin

end Behavioral;
